[your RTL code]
